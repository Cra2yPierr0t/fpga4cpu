module maindec(op, memtoreg, memwrite, branch, alusrc, regdes, regwrite, jump, aluop);

