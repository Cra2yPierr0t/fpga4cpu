module Fulladder(X,Y,Cin,out,Cout);


